some changes may be pushed to github