some changes may be pushed to github or may be not!